// https://veripool.org/guide/latest/example_cc.html#example-c-execution
module our;
     initial begin $display("Hello World"); $finish; end
  endmodule
