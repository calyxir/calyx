// Used by the comb-path.futil test
